module main

pub fn prob_1(a int, b int) int {
  return a + b
}
